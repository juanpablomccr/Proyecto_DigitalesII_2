`timescale 1ns/1ps
`include "modules/fsm/fsm.v"
module fsm_tb(
	clk,
	init,
	pause,
	continue,
	idle,
	emty_vc0,
	emty_vc1,
	emty_vc2,
	emty_vc3,
	stppd_vc0,
	stppd_vc1,
	stppd_vc2,
	stppd_vc3,
	cntn_vchanel0,
	cntn_vchanel1,
	cntn_vchanel2,
	cntn_vchanel3
	err_vchanel0,
	err_vchanel1,
	err_vchanel2,
	err_vchanel3
);



endmodule



module fsm_tester;

fsm fsm(


);

fms_tb(





);


endmodule
